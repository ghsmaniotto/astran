.SUBCKT NAND2X2 A B Z GND GND VDD VDD
MM64 n247 A GND GND NMOS l=0.06 w=0.2
MM65 Z A VDD VDD PMOS l=0.06 w=0.28
MM66 Z B VDD VDD PMOS l=0.06 w=0.28
MM67 Z B n247 GND NMOS l=0.06 w=0.2
.ENDS NAND2X2
